module top (
    
);



endmodule