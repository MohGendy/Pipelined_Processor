module adder (
    input  [7:0] a,
    output [7:0] sum
);
    assign sum = a + 1;
endmodule
